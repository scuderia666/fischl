module pkg

pub struct Package {
pub mut:
	name string [required]
	test string
}
