module pkg

pub struct Package {
	name string
}
